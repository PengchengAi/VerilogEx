module shift_reg(clk, rst_n, preset_n, D, Sin, Q, Sout);
  input clk, rst_n, preset_n;
  input [3:0] D;
  input Sin;
  output reg [3:0] Q;
  output reg Sout;
  
  always @(posedge clk or negedge rst_n)
  begin
  // -------- insert your code here ------------















  // -------------------------------------------
  end


endmodule