module adder(A, B, Cin, S, Cout);
  input A, B, Cin;
  output S, Cout;

// -------- insert your code here ------------



// -------------------------------------------

endmodule